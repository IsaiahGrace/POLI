/* 
 Isaiah Grace
 igrace@purdue.edu
 
 This module controls the orientation and status of the test structures
 */

// Includes
`include "POLI_types_pkg.vh"
`include "control_register_if.vh"

module control_register (
			 input logic CLK,
			 input logic nRST,
			 control_register_if crif
			 );
   // Import types
   import POLI_types_pkg::*;

   // local signals and registers
   
   // combinational logic

   // sequential logic
   
endmodule // control_register

     
